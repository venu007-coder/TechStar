Return-Path: eswari@jjcpl.net
Received: from mx12.stngva01.us.mxservers.net (204.202.242.5)
	by mail19j.g19.rapidsite.net (RS ver 1.0.95vs) with SMTP id 4-0997031784
	for <abhra@altechstar.com>; Tue, 17 May 2011 10:16:24 -0400 (EDT)
Received: from unknown [216.151.164.100] (EHLO mail.njtech.com)
	by va1-mx12.stngva01.us.mxservers.net (mxl_mta-3.1.0-05)
	with ESMTP id 83382dd4.1098300320.713089.00-011.va1-mx12.stngva01.us.mxservers.net (envelope-from <eswari@jjcpl.net>);
	Tue, 17 May 2011 10:16:24 -0400 (EDT)
Received: (qmail 28334 invoked from network); 17 May 2011 14:16:21 -0000
Received: from unknown (HELO NEW2-PC) ([122.164.92.161])
  by 10.97.0.64 with SMTP; 17 May 2011 14:16:17 -0000
From: "Eswari" <eswari@jjcpl.net> 
To: "abhra@altechstar.com" <abhra@altechstar.com>
Reply-To: eswari@jjcpl.net
Date: Tue, 17 May 2011 09:16:02 -0500
Subject: Oracle EB Tax module Consultant
MIME-Version: 1.0
Content-Type: multipart/related;
	type="multipart/alternative";
	boundary="=_reb-r518C6130-t4DD28338"
X-Mailer: aspNetEmail ver 3.6.0.66
Message-ID: <NEW2-PC037459f5fae641e38875828eb7d14217@NEW2-PC>
X-Processed-By: Rebuild v2.0-0
X-Spam: [F=0.2000000000; B=0.500(0); S=0.200(2010122901); MH=0.500(2011051716)]
X-MAIL-FROM: <eswari@jjcpl.net>
X-SOURCE-IP: [216.151.164.100]
X-SF-Loop: 1

This is a multi-part MIME message.

--=_reb-r518C6130-t4DD28338
Content-Type: multipart/alternative;
	boundary="=_reb-r4574D79C-t4DD28338"

This is a multi-part MIME message.

--=_reb-r4574D79C-t4DD28338
Content-Type: text/html;
	charset="iso-8859-1"
Content-Transfer-Encoding: quoted-printable

<!DOCTYPE HTML PUBLIC "-//W3C//DTD HTML 4.0 Transitional//EN">
<HTML xmlns:o=3D"urn:schemas-microsoft-com:office:office"><HEAD>

</HEAD>
<BODY>
<P class=3D"MsoNoSpacing" style=3D"MARGIN: 0in 0in 0pt"><FONT face=3D"Calib=
ri">Dear=20
abhra,<o:p></o:p></FONT></P>
<P class=3D"MsoNoSpacing" style=3D"MARGIN: 0in 0in 0pt"><o:p><FONT face=3D"=
Calibri">&nbsp;</FONT></o:p></P>
<P class=3D"MsoNoSpacing" style=3D"MARGIN: 0in 0in 0pt"><FONT face=3D"Calib=
ri">Good=20
Day!!!!!!<o:p></o:p></FONT></P>
<P class=3D"MsoNoSpacing" style=3D"MARGIN: 0in 0in 0pt"><o:p><FONT face=3D"=
Calibri">&nbsp;</FONT></o:p></P>
<P class=3D"MsoNoSpacing" style=3D"MARGIN: 0in 0in 0pt"><FONT face=3D"Calib=
ri">Hope you=20
are doing great!!!<o:p></o:p></FONT></P>
<P class=3D"MsoNoSpacing" style=3D"MARGIN: 0in 0in 0pt"><o:p><FONT face=3D"=
Calibri">&nbsp;</FONT></o:p></P>
<P class=3D"MsoNoSpacing" style=3D"MARGIN: 0in 0in 0pt"><FONT face=3D"Calib=
ri"><B>If you=20
have any consultant regarding for the below requirement please inform me th=
rough=20
phone or email</B>.<o:p></o:p></FONT></P>
<P class=3D"MsoNoSpacing" style=3D"MARGIN: 0in 0in 0pt"><o:p><FONT face=3D"=
Calibri">&nbsp;</FONT></o:p></P>
<P class=3D"MsoNoSpacing" style=3D"MARGIN: 0in 0in 0pt"><FONT face=3D"Calib=
ri">Position:=20
Oracle EB Tax module Consultant<o:p></o:p></FONT></P>
<P class=3D"MsoNoSpacing" style=3D"MARGIN: 0in 0in 0pt"><FONT face=3D"Calib=
ri">Duration:=20
Long term Contract<o:p></o:p></FONT></P>
<P class=3D"MsoNoSpacing" style=3D"MARGIN: 0in 0in 0pt"><FONT face=3D"Calib=
ri">Location:=20
NewYork City,<o:p></o:p></FONT></P>
<P class=3D"MsoNoSpacing" style=3D"MARGIN: 0in 0in 0pt"><FONT face=3D"Calib=
ri">Rate:=20
$75/hr.<o:p></o:p></FONT></P>
<P class=3D"MsoNormal" style=3D"MARGIN: 0in 0in 0pt"><B><SPAN style=3D"COLO=
R: black; FONT-SIZE: 14pt"><o:p><FONT face=3D"Calibri">&nbsp;</FONT></o:p><=
/SPAN></B></P>
<P class=3D"MsoNormal" style=3D"MARGIN: 0in 0in 0pt"><B><SPAN style=3D"FONT=
-SIZE: 14pt"><FONT face=3D"Calibri">In person interview mandatory after=20
phone<SPAN style=3D"COLOR: black"><o:p></o:p></SPAN></FONT></SPAN></B></P>
<P class=3D"MsoNoSpacing" style=3D"MARGIN: 0in 0in 0pt"><FONT face=3D"Calib=
ri"><B>Skills=20
needed</B> <o:p></o:p></FONT></P>
<P class=3D"MsoNoSpacing" style=3D"MARGIN: 0in 0in 0pt"><BR><FONT face=3D"C=
alibri">-=20
Skilled in Oracles EBTax module and the use of EBTax with both Oracle Accou=
nts=20
Receivable and Accounts Payables. <BR>- Ability to work with tax department=
 to=20
understand current tax rules and interpret those into EBTax rules. <BR>-=20
Experience in creating and testing EBTax rules related to Accounts Receivab=
le=20
and Accounts Payables. <BR>- Ability to recognize and solve tax issues that=
 are=20
found as testing is done. <o:p></o:p></FONT></P>
<P class=3D"MsoNoSpacing" style=3D"MARGIN: 0in 0in 0pt"><o:p><FONT face=3D"=
Calibri">&nbsp;</FONT></o:p></P>
<P class=3D"MsoNoSpacing" style=3D"MARGIN: 0in 0in 0pt"><FONT face=3D"Calib=
ri"><B>Responsibilities of the role:</B> <o:p></o:p></FONT></P>
<P class=3D"MsoNoSpacing" style=3D"MARGIN: 0in 0in 0pt"><BR><FONT face=3D"C=
alibri">- Need=20
to work with tax department to have key decision made examples include dire=
ction=20
around tax determination factors, criteria for tax applicability and what i=
s=20
taxable in the following scenarios: direct pay permit , p-card transactions=
,=20
incoming AP invoices from feeder systems, AR transaction types, and one-tim=
e=20
delivery addresses. <BR>- Complete the mapping of tax requirements based on=
 the=20
identified drivers. Then determine how to complete in Oracle the tax rules =
that=20
will need to be implemented. <BR>- Then configure in Oracle and test the ru=
les=20
to validate that the configuration matches all the requirements.=20
<o:p></o:p></FONT></P>
<P class=3D"MsoNoSpacing" style=3D"MARGIN: 0in 0in 0pt"><SPAN style=3D"COLO=
R: black"><o:p><FONT face=3D"Calibri">&nbsp;</FONT></o:p></SPAN></P>
<P class=3D"MsoNoSpacing" style=3D"MARGIN: 0in 0in 0pt"><FONT face=3D"Calib=
ri"><B>Note=20
</B>:-If you are interested and have above skills kindly fill the submissio=
n=20
form attached with this email along with your updated resume and send back =
me=20
immediately.<B><SPAN style=3D"COLOR: black"><o:p></o:p></SPAN></B></FONT></=
P>
<P class=3D"MsoNoSpacing" style=3D"MARGIN: 0in 0in 0pt"><SPAN style=3D"COLO=
R: black"><FONT face=3D"Calibri">&nbsp;</FONT></SPAN><o:p></o:p></P>
<P>
<P class=3D"MsoNormal" style=3D"MARGIN: 0in 0in 0pt"><SPAN style=3D"mso-far=
east-font-family: 'Times New Roman'; mso-fareast-theme-font: minor-fareast;=
 mso-no-proof: yes"><FONT face=3D"Calibri">Thanks for choosing JJCPL<o:p></=
o:p></FONT></SPAN></P>
<P class=3D"MsoNormal" style=3D"MARGIN: 0in 0in 0pt"><SPAN style=3D"mso-far=
east-font-family: 'Times New Roman'; mso-fareast-theme-font: minor-fareast;=
 mso-no-proof: yes"><FONT face=3D"Calibri">Regards </FONT></SPAN></P>
<P class=3D"MsoNormal" style=3D"MARGIN: 0in 0in 0pt"><B><I><SPAN style=3D"F=
ONT-FAMILY: 'Century Gothic','sans-serif'; COLOR: #215868; FONT-SIZE: 12pt;=
 mso-fareast-font-family: 'Times New Roman'; mso-fareast-theme-font: minor-=
fareast; mso-no-proof: yes">Eswari</SPAN></I></B></P>
<P class=3D"MsoNormal" style=3D"MARGIN: 0in 0in 0pt"><SPAN style=3D"FONT-FA=
MILY: 'Century Gothic','sans-serif'; COLOR: #215868; FONT-SIZE: 12pt; mso-f=
areast-font-family: 'Times New Roman'; mso-fareast-theme-font: minor-fareas=
t; mso-no-proof: yes"><FONT face=3D"Calibri" color=3D"#000000">Recruiter</F=
ONT></SPAN></P>
<P class=3D"MsoNormal" style=3D"MARGIN: 0in 0in 0pt"><SPAN style=3D"COLOR: =
red; mso-fareast-font-family: 'Times New Roman'; mso-fareast-theme-font: mi=
nor-fareast; mso-no-proof: yes"><FONT face=3D"Calibri"><IMG height=3D"35" w=
idth=3D"138" src=3D"cid:image_0000" alt=3D""></FONT></SPAN></P></P><SPAN st=
yle=3D"COLOR: red; mso-fareast-font-family: 'Times New Roman'; mso-fareast-=
theme-font: minor-fareast; mso-no-proof: yes"><FONT face=3D"Calibri">
<P class=3D"MsoNormal" style=3D"MARGIN: 0in 0in 0pt"><B><SPAN style=3D"FONT=
-FAMILY: 'Tahoma','sans-serif'; COLOR: #f2f2f2; FONT-SIZE: 7pt; mso-fareast=
-font-family: 'Times New Roman'; mso-fareast-theme-font: minor-fareast; mso=
-no-proof: yes"></SPAN></B><SPAN style=3D"COLOR: red; mso-fareast-font-fami=
ly: 'Times New Roman'; mso-fareast-theme-font: minor-fareast; mso-no-proof:=
 yes"><FONT face=3D"Calibri">&#8220;<I style=3D"mso-bidi-font-style: normal=
">we forecast you</I>&#8221;=20
</FONT></SPAN></P>
<P class=3D"MsoNormal" style=3D"MARGIN: 0in 0in 0pt"></FONT></SPAN><SPAN st=
yle=3D"FONT-FAMILY: 'Bookman Old Style','serif'; FONT-SIZE: 9pt; mso-fareas=
t-font-family: 'Times New Roman'; mso-fareast-theme-font: minor-fareast; ms=
o-no-proof: yes"><o:p></o:p></SPAN></P>
<P class=3D"MsoNormal" style=3D"MARGIN: 0in 0in 0pt"><SPAN style=3D"mso-far=
east-font-family: 'Times New Roman'; mso-fareast-theme-font: minor-fareast;=
 mso-no-proof: yes"><FONT face=3D"Microsoft Sans Serif" size=3D"2">469 327 =
3112</FONT></SPAN></P>
<P class=3D"MsoNormal" style=3D"MARGIN: 0in 0in 0pt"><SPAN style=3D"mso-far=
east-font-family: 'Times New Roman'; mso-fareast-theme-font: minor-fareast;=
 mso-no-proof: yes"><A href=3D"http://www.jjcpl.net/"><SPAN style=3D"COLOR:=
 blue"><FONT face=3D"Calibri">http://www.jjcpl.net</FONT></SPAN></A><FONT f=
ace=3D"Calibri">=20
<o:p></o:p></FONT></SPAN></P>
<P class=3D"MsoNormal" style=3D"MARGIN: 0in 0in 0pt"><SPAN style=3D"mso-far=
east-font-family: 'Times New Roman'; mso-fareast-theme-font: minor-fareast;=
 mso-no-proof: yes"><FONT face=3D"Calibri">Skype: jjcpl.rpo</FONT></SPAN></=
P>
<P class=3D"MsoNormal" style=3D"MARGIN: 0in 0in 0pt"><SPAN style=3D"mso-far=
east-font-family: 'Times New Roman'; mso-fareast-theme-font: minor-fareast;=
 mso-no-proof: yes"><FONT face=3D"Calibri">Gtalk : jjcpl.rpo</FONT></SPAN><=
/P><SPAN style=3D"mso-fareast-font-family: 'Times New Roman'; mso-fareast-t=
heme-font: minor-fareast; mso-no-proof: yes">
<P class=3D"MsoNormal" style=3D"MARGIN: 0in 0in 0pt"><B><SPAN style=3D"COLO=
R: #31849b; FONT-SIZE: 11pt"><FONT face=3D"Times New Roman" color=3D"#0000f=
f"><A href=3D"http://jjcplrpo.blogspot.com/">http://jjcplrpo.blogspot.com</=
A>=20
</FONT></SPAN></B></P></SPAN><SPAN style=3D"mso-fareast-font-family: 'Times=
 New Roman'; mso-fareast-theme-font: minor-fareast; mso-no-proof: yes">
<P class=3D"yiv1141086511msonormal" style=3D"MARGIN: 0in 0in 0pt"><STRONG><=
SPAN style=3D"FONT-FAMILY: 'Calibri','sans-serif'; COLOR: gray">Note: We re=
spect your=20
online privacy. This is not an unsolicited e-mail. If you are not intereste=
d in=20
receiving our e-mails then please reply with a</SPAN></STRONG><SPAN style=
=3D"FONT-FAMILY: 'Calibri','sans-serif'; COLOR: gray; FONT-SIZE: 10pt">=20
</SPAN><STRONG><SPAN style=3D"FONT-FAMILY: 'Calibri','sans-serif'; COLOR: r=
ed">"REMOVE"</SPAN></STRONG><SPAN style=3D"FONT-FAMILY: 'Calibri','sans-ser=
if'; COLOR: gray; FONT-SIZE: 10pt">=20
</SPAN><STRONG><SPAN style=3D"FONT-FAMILY: 'Calibri','sans-serif'; COLOR: g=
ray">in=20
the subject line. All removal requests will be honored ASAP. We sincerely=
=20
apologize for any inconvenience caused to you</SPAN></STRONG><SPAN style=3D=
"FONT-FAMILY: 'Calibri','sans-serif'; FONT-SIZE: 10pt"><o:p></o:p></SPAN></=
P></SPAN></BODY></HTML>


--=_reb-r4574D79C-t4DD28338--


--=_reb-r518C6130-t4DD28338
Content-Type: image/jpeg; name="logo%20new%201.jpg"
Content-Transfer-Encoding: base64
Content-ID: <image_0000>
Content-Disposition: inline

/9j/4AAQSkZJRgABAAEASABIAAD//gAfTEVBRCBUZWNobm9sb2dpZXMgSW5jLiBWMS4wMQD/
2wCEAAUFBQgFCAwHBwwMCQkJDA0MDAwMDQ0NDQ0NDQ0NDQ0NDQ0NDQ0NDQ0NDQ0NDQ0NDQ0N
DQ0NDQ0NDQ0NDQ0NDQ0BBQgICgcKDAcHDA0MCgwNDQ0NDQ0NDQ0NDQ0NDQ0NDQ0NDQ0NDQ0N
DQ0NDQ0NDQ0NDQ0NDQ0NDQ0NDQ0NDQ0NDf/EAaIAAAEFAQEBAQEBAAAAAAAAAAABAgMEBQYH
CAkKCwEAAwEBAQEBAQEBAQAAAAAAAAECAwQFBgcICQoLEAACAQMDAgQDBQUEBAAAAX0BAgMA
BBEFEiExQQYTUWEHInEUMoGRoQgjQrHBFVLR8CQzYnKCCQoWFxgZGiUmJygpKjQ1Njc4OTpD
REVGR0hJSlNUVVZXWFlaY2RlZmdoaWpzdHV2d3h5eoOEhYaHiImKkpOUlZaXmJmaoqOkpaan
qKmqsrO0tba3uLm6wsPExcbHyMnK0tPU1dbX2Nna4eLj5OXm5+jp6vHy8/T19vf4+foRAAIB
AgQEAwQHBQQEAAECdwABAgMRBAUhMQYSQVEHYXETIjKBCBRCkaGxwQkjM1LwFWJy0QoWJDTh
JfEXGBkaJicoKSo1Njc4OTpDREVGR0hJSlNUVVZXWFlaY2RlZmdoaWpzdHV2d3h5eoKDhIWG
h4iJipKTlJWWl5iZmqKjpKWmp6ipqrKztLW2t7i5usLDxMXGx8jJytLT1NXW19jZ2uLj5OXm
5+jp6vLz9PX29/j5+v/AABEIAFgBGAMBEQACEQEDEQH/2gAMAwEAAhEDEQA/APsugAoAQnHJ
4xQBgyeIInYx2Mcl86kg+SB5SkdmmYrF9QrMw7rXQqLWtRqC/vb/APgK1++3qc7qramnJ+Wy
/wC3tF+ZGLvU2LbktLZUXcVeV3ZV5+ZtqooXg85xweeDVctNbOb9EkvldsL1O0Y9dW21+RXt
dWuL1iltcafMyjcVRnJx/e4c/L/tYxTlTjDWUaiXnb/IlTlLSMoP0v8A5kkWq6go3tbxXUWf
v2k4Y49kkCA/g9J06eyk4vtONvxV/wAhqc1q4qS7wl+jt+Zp2WsW18xiRjHMoy0MqmOVR67G
AJH+0u5PRjWUqcoav4eklqvvX5PU0jUjLRaPs9H9z/PY1KyNQoAKACgAoAKACgAoAKACgAoA
KACgAoAKACgAoAKACgAoAKACgAoAKACgAoAKACgCne30WnRebMSBkKqqCzO54VEUcs7HgAfy
yauMHN8sf8kl1bfRESkoK7+S6t9l5mQunTat+81P5YicraKfkA7eew/1reqD90OmH61tzqlp
R3/n6/8Abq6eu/oZcjqa1dukOn/b3f029SvrV6lhNaR20ipJHNGrWqkAyQTbouIxyRGf3i4G
B5Z7ZqqcXJTclo4u0n0ktd/Pb5inJQcVF2aa91dU9NvLf5GHrED6lNNJOosFNt5LNcvGI5Xi
uFliA2uS0TL5gckL8sgG0nIG9NqmoqPvvmuuVO6Ti0+m+1vTcxmuZtv3Pdt7zVm1K667PW/q
MvNbj1SN0B06OUW80cRF3DJL5kqbAImG0IgBJck5bAG0YzTjSdNp/vGuaLfuNKyd9Vrd9vzE
6immvcT5Wl76bu1bTsu42XTH0CCPUY3tttooANvH5T3LMvlRQylXMZRpGUlipYYBBXk0Kaqt
02pe8/tO6jrdyWl7pX0Bx9klNOPu/wAqtzdEnra1zs10pby0ih1HFxNGilpQNjCTA3PGy4MZ
z0KEccetcXtOSTdL3U29N1bs77/M6uRSilU1a67a91bb5FUXU+iNtvWM1oSAtyR88WTgLcAA
AqegnAAB/wBYAPnrTljV/hq0/wCXo/8AD5/3fu7EXdLSbvHpLqv8X/yX39zoxzyK5TpCgAoA
KACgAoAKACgAoAKACgAoAKACgAoAKACgAoAKACgAoAKACgAoAKACgCOSRYUMjkKiAsxPAAAy
SfYCmld2W/QTfKrvZGDpkDX8v9q3IIyCLWM/8soj/GR/z1mHLHqqERjHz56JtU17GH/bz7vt
6R/F69jCC537WX/bq7Lv6v8ALTubN3eQ2ETXFwwjjQZJP8vcnoAOSeBWEYubUYq7ZtKSguZ6
JHlmqeIr3Urho4MWEcajaxANy6v2zhjHk4AhjV52JB27SGr14UYU4py99t7fZVvLr/idorv0
PNnUlOVo+4lt/M7/AJeiu/zOEv8AwQ2qSktmZ3cRYldi5lwcor5fayrl5h86wqDuYyEovoQx
Ps1ZaJK+iVrd7aekdubtbV8csPzvXVt21b37X19X29dBk/hIXFtFFLGJLW1TzIleYlFgErQG
RQsQbA+STJOQhPXpSjX5JNxdpN2do681ua29u69QdHmilJXitVeWiV2r7ej9DY03wxJo24Qu
0ZJETxKcRqxHyxujkxP5gOY3kURzqV2ujfKcZ1lVtzK/VPq/NNaq3VJ3j1T3NY0XT+F26W6e
lno79G9H5Hd+GdfFlmwulCRxvsWZdwTeeWjZGJ8opwGVSFQkApGuCfPrUub95B6tX5etu91v
f8e7OylU5fcktE9H0v2t0t/SR6IyrIpVgGVhgg8gg9QR0IIrzdtVozv8jn7EHRrgaexJtpcm
0JOShAy9uSeSFHzQ552Bk52CumX72PtV8S+Pz7S+e0vPXqc0f3cvZ/Zfw+XeP6ry06HR1zHS
FABQAUAFABQAUAFABQAUAFABQAUAFABQAUAFABQAUAFABQAUAFABQAUAYWqj7ZLFp38MpMkw
/wCmMZBKH2lkKIfVPMFdFP3FKr1Wkf8AE+vyV362MJ+81T6PV+i6fN2Xpc3CQoz0ArnNzyPV
9Rk1O7F/IWTTLPdkopYxBsBLrb/FNJhlhXa3kQus5Xc6kezTgqcfZr+LLvpfvC/SK3ltzSXL
eyZ5c5Ocud6U4/h/et3fTsnzdTUXTk1BIY0VPMuAWi2tuFlBxvlVwSTdS5CmXduMjYB2I+ce
dwbbvaO99OeXRW/kXba3m0a8qlZLd7f3I9Xf+Z9+/kmVzp7WcF1fWdxLFBYxy29orBJRkcSu
C4LZeYBA27cRGWyd5FVzqThTnFOU2pTeq9Fp2jr8/Inl5VKcJNKKcY7P1evd6fLzLcekXdrc
Wlo9yNj2csGPIj+6oiJQ5JByAeo9fU1DqRcZzUdVNS+J9b6lqEouMebTla+FeRTTSHS3eW4k
lu309mtbmEkKs1omGXKIAWYQsky5Jy29B941ftFzJRSiprmi/wCWb83tqnF/JkqFldty5fdk
trx+XlZ/eTXsFtpqrA7J5MsYNmx5FxGBn7I4UFnkUHNtKoMmD1Yq4kmLlP3kndP3/wC6/wCd
dl/Mtvws5KMfd6Ne75r+X1/la1/G97wjqc0O3Tb0tlxI9sX++ERyHtZSAB59sCgbHDKQykgZ
rOvBP95T8lK212tJr+7LX576l0ZNfu5+bjfe38r84nW6pZm9t2jQ7ZVw8Tf3JUO5G+m4AMO6
ll6E1y05ckk3ts13T3/rudE480bLR7rya2JdPuxfW8dwBt3rkr/dYcMp91YFT7ipnHkk49vy
6P5rUcZcyUu/9M4r4lS6rY6NPqWjXjWE1hE8zDyYJUmVQCVbzo5CpChthTHzH5wRgjagouah
ON1J23at9zMq3NGDlCVmlfZO/wB55nrfjvXp9I8N/YLhLS916VIZ5/JikAYtHFuEboyAFpN7
BVB4wpA4rshRpqdXmV401dK7Xd9/I5ZVZuNLldnN2bsvQ9KvPDXiFbZ/smu3JughKeZaad5T
SAcBgtoGCseOHJUHPzY541Ondc1NW8pTv/6UdThNL3ajv00jb8jjfHPiXxHpzeHdLtp006/1
hhHeyCKGYRyqtqsgRXWSMqrzSEbfvbVAcLknopQpv2s2uaMPhV2tNbduiRhUnUj7OCfLKXxa
J66f5nqt/pmoTab9ktL6SC+VABeGG3dmdR954TH5O1z94Ii4H3Cp5riUoqV5RvH+W7X43udb
jLl5VK0u9l+Wx5t8N/H9xf8AhOfX9fkErWMk4eRURGdI1R1GxAibyX2KFVQTtzzknrr0VGqq
VJWvay7XOWjVbpOpU6X8i14Yk8TeNLJdamvv7Ghusva2lvbQTFYskRyTS3KSM5kA3YjEYKlW
BXdsWansqL9mo87W7ba18krW/H9Soe0qrncuRPZJJ6ebZf8ABvi++n1W88La8I/7SsFEsc8S
lI7q2bbiUISQjgOm9VJXLMBjY2Zq04qEa1K/LLSz3i+xVOo+Z0qnxLVNdV3Mj4Z6/q3iC+1K
PWLx/tGmXckDWSQ26QCNiRE6uIRcN8ySBczEEBWYndWleEKcYezjpKKfNd3v1627dCKMpTcl
N6xduWyt5dL9+p03i+51G1v9Nj027kie8u44WtRFbvE8Me+a6mdnhaZSsClBslQbjHgAlica
ai4z5orRN3u077RW9t/I1qOSlFRdru1rK1lq3tfbzOJ8Z/Ei/wDD/ia0t4QBosM0NrqEhRCP
tF0jSKu8/Mphh2T/ACEA5YPn5RXRSoRnTk38bTcV5L/N6GFSs4VEl8CaUvV/5LU9C+Imt3Ph
zw9e6lYkLcW8QMbMAwVnkSPdtIIJXdkBgRkDIIyK5aMFUqRhLZv9LnRVk6cJSjuloRfD7+1L
nRbe+1e9a+uL+CK4B8mCJYVljDqiiKNNxAYbi+7LA4wvBdblU3GEeVRbW7d7PzYUuZwUpyu2
k9krX9Ecf4S17W4PGV/4Y1O8/tG1t7MXMMjQQQyKS1vgHyI4weJ2VsgglVZQmStb1IQ9jGtC
PK3Kz1b7935GFOU1VlSlK6UbrRLt29T2quA7jxK31zXNH8dReHbu9+3afe2klzGrwQRvF/rs
LvhijLFWgYZJIKMMjcM16DhCVB1Yx5ZRlbdtPbu/M4VKcaypuV4tXWiVt+y8jJ8Wah4o0/xZ
Y6HZau0Vnq2+Rc2lmzwKhdnjUmD5wEUCNmO7J+fOMtdONJ0pVJQ96H96ST89yJupGpGEZ2Uv
KOn4G74817WNO1fQ9B068NqNRaRbi58mCSV/LEYyFkjaJS2WJ2oAGIwNo2nOjCEoVKko35dl
dpLfs7mlWUoyhTjK3Nu7Jvp5WGeNNR8QfD20XW1v/wC1bSKWNLi2ure2icpIwXdFLaxQ4cMQ
MOrDndztKkpRp137Pl5XZ2abf3ptiqOdFc/NzJPVNJfc0kV/FvifWLzxLpGg6Hef2db6nbNc
vL5EMrlQssmNsyOAfLhIUDHzN8xIAp06cI051KkeZxdkrtdl0fmKc5OpCnTfKpK97J9319Dp
da0HxRaWrz6Rq811dxYdLe5ttPEU+CCYi8dtC0ZcZAfeMHqVzuGUZ0m7Tgku6crrz3ZrKNRK
8JttdGo2flsvzMDxbr2tzeMbDwxpV5/Z1tcWZuZpFggmkJDXGQPOjkAOIFC4wBuZjuwFrSnC
CoyrTjzNSsldrt2a7mdSU/axpQlypq70T79/Q7Lx9/adpolxe6TetZXFhby3JbyYJRMIYy7I
6yxuF3BThkC4YjOVypwo8rmozjdSaW7VrvyZvV5lByhKzim9k729ST4d63c+IvD1lqV8Q1zP
GxkZVChmSR03bRgAsFBIUBck4AGBSrQVOpKEdk9PuCjJzhGUt2blohe/uZm/gEMK/wC6E8w4
/wCBSfpRLSEEv7zf32/QcV78n2sl91/1K/ii4Nvp0oG4GYeUNn3v3nynb6HbnB9cU6Eb1F5a
6+QqrtBpddPvOZ0CPy5E0y7/AHb6agmnyci4nIGyVWwN8cSYbHBV2jBAMYz1VXo6sNpu0f7s
eq8m396v3MKas1Tlo4av+8+/mkvxt2FbTo4bK41qISWtzcZeMQMY/lPyW6Mg+RiSRI+VOXdz
3o525xoO0ox0fNr5yd9/JeSQcqUZVVdSe1tP8Om3n82Pv9GvbDT4bGO53o8lvCVeFT1kUsSy
FCRkEknkjOT3pQqQlOU3GzSk9JNdH0dwlCUIKClpeK1Xn5WL+ow6it7ZsZbfO+ZQRBJxuhY8
5nPXbxyOfXpWcHT5JpKWy+0v5l/dNJKfNHWO76Ps/MYum3i6k0ct06rdQh2MMaR5aFtuNxDk
Eo685yQvtT54ezTUFeMrK7b0evl1X4i5ZKdnLdX0SW339yDT/D1vD9osEBW4tmV7a4cs7ojZ
eHazEkCNw8TKmA0ahW+8ac6sny1H8LupRWib2ei7qz16ijTS5oLdaxe7S6fc9PQyb+5e9ngu
rRTG8biW5+UlY7qBGBgVu7zRiSKQgEBVjJOSudYxUFKE3dNWjrvGT+L0i7Ned/Mzk+ZqUVaz
u/KSvp81dP5HqSMHAZehGR9DzXl7aHoGXpUJtjcR9FFw7IPQOqSHH/Anb8a2qO/K/wC6r/Jt
fkkZQXLzLpzO3zSf6s5/4k/8ixqn/XlP/wCizVUP4sP8S/Mmt/Dn/hZ856t9o/sfwT9i8v7T
9pXyfN3eX5vnW/l+Zt+bZvxv2/NtzjmvUjbnxHNe1tbb2s9vkebK/JQ5d76X73R9LaN/wkn2
j/ib/wBm/Ztp/wCPX7T5u7jb/rfk29c9+mK8mXs7e5zX87W/A9OPtL+/y28r3/E8o+Mn2r+3
/DH2Dy/tP2u48rzt3lb99ljzNnz7P7235sdOa7cNb2dbmvblV7b/AGjkxF+ely73dr7bxPQH
/wCE22nb/Ym7Bx/x+9e1c37n/p5/5KdH77+5/wCTHzno3mf8Ko1Hyun25d+M52edZ5xj3xn/
AGc5r1JW+tRv/L+kjzo/7tK3836xPrLwv5X9j2P2fHlfY7by8dNnkptxnttxivFqX55X35n+
Z60LckbbWX5HlOq7f+Fn6f5Wd39kyebjGMbrrbuxznO3O7t5eK7Y/wC7Sv8Azq3/AJKckv8A
eI2/k1/Eg1b/AIoz4g2t+Pks/EkBtZfQXMexUOBgAsRbqCeT5kp7mnH97h3H7VN3Xo/6f3IU
v3VdS6TVn6/1b72dgt7Dca5qGt3JxZeH7VrVX6gSuq3V845xlI1t4j3yHGaws1CNNfFN3+S0
j+N2bXTnKb+GCt895fojyPUNS0LXfBd1b3d/ZDVdQaXVGjM6bkunfzY4QCchlhVLTB6cjgdO
2MZwrRcYy5I2ht02v9/vHI3CVJpyjzO8t+u9vu0NzU/Ef/CUfC+a9c7pkt44J/XzYZ4kYn3c
BZP+B1nGHssSora7a9Gn/wAMW58+Hcutkn6pr+vmdJ4M/wCEv/sLTvs39j+R9htfK8z7Z5nl
eSnl+Zt+Xfs279vy7s44rKr7LnlfnvzO9uXe7ua0/a8kbcluVW+La2hzXg3+0P8AhZOpf2t9
n+1f2Uu77L5nlbd9jt2+b8+duN2f4s44xWtXl+rQ5L25+u/2uxlT5vby57X5Om32e59F15Z6
R4RrP/JUtM/7BL/+hX9ejH/dZ/41/wC2nBL/AHiP+D/5IXxr/wAlA8Pf9c7n/wBAlopfwKvy
/NBU/jU/n+pk/GCW+t/EugS6UiTXiG5aGOQkI7jyjsJBUjcMgcjkjJxmrwyj7Oqp6R0vbpuR
iLqpT5N9bL7hujT6h8bbL7NqlxbWFpaXI+22NtFKLpihJRJHlkIjRiCQVRvnRgfmQhSSjg5X
gnJte7JtW17W3/4IR5sUrSaST96KTv8Aix3jeO8h+IGiR6MLdblLGZYhcbxAFCXYcMIvn4i3
BNv8W3PGaKVvq9TnvbmV7b/Z7+YVLqtBQtfldr7de3ke0aF/bu9/7a+wbMDy/sfn7t2Tnf53
GMYxt5z1rgn7P/l3zf8Ab1v0O2PP9vl8rX/U8Y8Zf2h/wsnTf7J+z/av7KO37V5nk7d99v3e
V8+duduP4sZ4zXfS5fq0+e9ufpv9nucVTm9vHktfl67fa7HS+M/+Ev8A7C1H7R/Y/kfYbrzf
L+2eZ5Xkv5nl7vl8zZu2bvl3YzxmsqXseeFue/MrfDa91Y1qe15JX5Lcrv8AFtbWxt/B3/kU
dO/65Sf+j5azxP8AFl6r8kXh/wCFH0f5s6pdbc6sdJ+zTBFh837Vj9yTkDy8/wB7nuR6Y6E+
Z7R+09lyu1r83T0PofqcVglj/bU+Z1OT2N/3ltfft2/ruTa9eS2FvHNCQGN3ZRHIBBSe7ggc
c9DslYqRghgD0yDVSThFOP8ANBfKU4xf4MywVKFepOnUV0qGJmrO1pUsPVqwf/gUFdPdX62Z
z9jqd69rp9zJ5rvevFvjK2obBtJp3MRBCqjsij943mBEYD5iCeeM58tOTveTjde7/LKTt0tf
u728z1q2Gw8a2LowVOMcPGpyzvXaTWIpUY8905OcYyfwR5HKSv7qZRt/EV9Nb3kzMIzp0VzM
FZUzL5V7fwpHKRlVCx2aK7QkEvIWBAChoVWbjOV7cik+mtp1I2fygr26v7+qeAw8KuHpRi5L
EzoU7py/d+0w2EqynTTs23PEycVUVlGCi0221el1y6UyWoYrdxzyADy9+IpVU258tFLv5YmR
n2HLm2uPmABAt1JK8ftKT6X0fw6LV25le2/LLU5o4Ki1Cva9CVODvz8v7yDarLnk1GPO6Uox
5l7vtqPuttN0LrxTePY3N7Ajh7fSxcFQse2G6U3ayrKJWWQhJLYxlUBOBJkbihrN1pckpxTv
GnzdNJe/e93fRxtZefWx108soRxFHDVZRcamN9im3O9Sg1QdN03BSgnOFZT5pNK7hry819vx
Rqlzpe02zBc297Jyob54YPNjPI7MMEdCCe+CN605Q+F/Zm/nGN0eXluGpYq6rRbtWw0dG17t
WryTWndPR9Gu10ZD+ILxLiWBGJeFC/zpGImjSxhmdgeJGnE8qEquUEbrlQDuGPtZJuKeqV9U
rWUE3583M15WfzPQjgKDp06sopRnJR92U3UU5YqpTimtYKk6VOVpStJzi7Sez1Y768ie1U+f
J9oSR3jItBICqKQQVZYwmXyBuL5AzkEitlKacfid07r3b6JfK2vqcMqNCUa7Xso+ylCMZJ4j
kfNKV000581o2bso2btrZmpoF/LfaXb3kw3SyQK7BQBliuTgZ2gn64z7VpSk5U4ze7imcGNo
Qw+Lq4alpCFSUY3bdlfTXfT7xPDusvrtp9qkt5bJt7p5cww2FON3QcN2/rRSqOrHmcXHVqz3
0Hj8JHAVvq8K0Ky5Yy56esfe+zvuupgfE+4S28L6kXON9q8S+peXEcaj1LOygAcnPFd9BXqw
t3v92p4dZ2py9LfeeV6t4H15dF8Mvp9stzeaHJHcTWzSxxHOYpgpaVkX5Wj8t8NuBOVBAJrt
jVp89ZSdozuk7X7rp96OSVKahS5Vdw1avbs+tj0688S+ITbP9k0K5F0UITzLvTvKVyOCxW7L
FVPPCAsBj5c5HGoU7q9RW8ozv/6SdbnO3u03f1jb8/0ON8c+GvEeoN4d1S2gTUL/AEZhJexi
WGESSstq0hRnaOMKzwyAbfu7lIQrkV0Up04+1g3yxn8Ojdlrbu+qMKkKj9nJK8o/Erpa6f5H
qt/qWoQab9rtLGSe+ZARZma3Rldh915TJ5O1D94o7ZH3Ax4riUY83LKVo/zWf5WudbclG6je
Xa6X43sebfDfwBc6f4Tn8P6/GImvZJy8aujsiSKiKdyF03gpvUqzAHbnnIHXXrJ1VVpP4bW6
banLRpONJ06ite+na5a8Mx+JvBVkuiy2P9sw2gKWt3b3NvCWiySkc0Vy8bIYwduYzINoVQG2
7mU/ZVX7RS5G9003r5NfrYqHtKS9m48yWzTS080/0uX/AAb4QvrfVbzxTrxjGpX6iKOCFi8d
rbLtxEHIAdyETeygLkMRne1RVqRcI0aV+WOt3o2+/kVTptSdWp8T0SXRdv6/Uk+K3hG48XaK
YtOH/Ews5o7m1+YITIhwyh2ICkozFSSF3qmSMZBh6ipT974Wmn/wwV6bqQtH4k7roZN34W1O
18Kw6WsTX15dXEU2qqkkKSTCWf7RehHlaOIsx/cjLKpiOAMYFWqkXVc78sUmoaOysrR0V35+
pDhJU1C122nLZXu7y308vQ9RS6mFn9o+zSLMI9wtd0PmBgMiLeJPI3Z+Xd5vl992K47K9r6X
31t67X/A67u17a9tPu3t+J892Pw/1w6P4i05LUWUGqSrPp9rJNAzq3mb5FLQyPEgZVjjXdJx
tGSBlq9R1oc9Kd7uKtJpP9de55ypT5KkUrKTvFXX6aHrfw+GqWui29hq9k1jcWEEVuB50Eqz
LFGEV0MUj7SQo3B9uGJxlea4a3K5uVOV1Jt7NWu/NI7KXMoKM42cUlune3ozj/CWg63N4yv/
ABNqdn/Z1rcWYtoY2ngmkJDW+CfIkkA4gZmyQAWVVL4LVvUnBUY0YS5mpXejXfv6mFOM/ayq
yjypqyV0+3Z+R7VXAdx4ncWcmp/EuG6txui0rSgly3ZJJmufLjJ7O6zK6qcEoGboOfQTUcM4
veU9Pla/5HC1zYhNbRjr87/5mR4s07xRf+LLHW7LSGks9J3xrm7s0edXLq8igz/ICjAxqw3Z
Hz4zhbpulGlKnKdpS/uy08tiJqo6kZxhpHzjr+PY2fiFoOt6hquia9pNn9qbTXd57ZpoYnUP
5RK73kWMnAddyM4DgHDKc1nRnCMKlKcrc2zs338r/kXVhNyhUhG/LurpdvMra54Q1fTNZg8Y
+GLfbdXKqup6Y8sUfmhgC+JN/keYMDcwcr5qLKu/MgZwqQlB0Kz0XwSSeny3/wCBoKVOUZKt
SWr+KN1r+Nv+Dr3DxVo2vzeJNI8Vadp5uBaW0kdxatcW0ckZkEyMC7TeUx2zEqY3ddy/NgHk
pypqnOjKVru6dnZ7dLX6BOM/aQqxjey1V0mr387dTp9a17xRdWrwaRpE1rdy4RLi5udPMUG4
gGUpHczM5QZITYcnqGxtOUYUk7zmml0Sld+Wy3NZSqNWhBp9242XnuzA8XaDrcPjGw8T6VZ/
2jbW9mbaaNZ4IZAS1xkjzpIweJ1K4yDtZTtyGrSnOHsZUZy5W5XWja6dl5GdSM1VjVhG6Ss1
dLv39TsvH/8Aad1olxZaTZNe3F/BLbFfOgiEImjKM7tLIgbaGOFQtlgOQuWrCjyxmpTlyqLT
2bvZ30sjerzODjCN201ula/qyT4daJc+HPD1lpl8AlzbxsJFVgwVnkd9u4ZBKhgCVJGQcEjk
qtJTqSlHZvT7gpRdOEYy3X+Z0lvds91PbOAPKEbJjOSjqck/R1YcY6fjUOKUYyXW6fk0/wDK
xal70ovpa3o/+DczvFEsttYtcQxLctbyRS+U5IDeXIrAgggBkIEibvl3oufUOnThVkqdR2XR
9mtY/iv13NPbVMOpVKOkuWUX/hmnCaT6c0W4vybXVmPpdxp9ylg1lBaBbnl9kKL5UkELMoVQ
BseJ2YKG5RSwXG4kt4aFLnTilycvKrJdbJ7dm7NdzR4/EVuVyr1Jc6mpXqTd+ZJzTu/tOMeZ
P4rK97IbJFcWV3FZ/Y7K8jVJZk8pFgkTEsZyqSbowxeQuxEil3+f5SOWqNCUOZLks0kmlJJu
7eyT3V9t++5LxeKjNr2s5c8feaqTTkopQSld6pR91Jv4dNEPudcWK+hE1hMjyBy7m3Esn7lW
8vY8LSZ2GV+52iRsY3nNrDxalNSg2uWzul33uk9Lu3q+5l9ZqQSop1FD3rxTfL73LzaJ297k
hzd+WN9kV77U9NiCIlizC4kEMqvYP80cjNI648sBt0nzlTkM5LEFjmojhIvmuqfwvrDXW9n5
X1fnqbvMK8XBxq1k4yi4+9UTi1Hki466SjBKKa1UVyrTQl1rVRcRiQadNcbSIj9pjRI9k7xo
4KyuudwwMlGxyCMFgWsPCbtVlDaXXm6a6JNdDOGLrYdP6u5wvKErp8jvFvlaldSVnK6s97Pd
Jjrm2nt9lxNaWEEXmwRmMR+bJgnyF/ebYkQpG+xQEkAQlAwUkGY0aDvFK7s2naKXuxdtNW9N
N1oaPGYpaurNK+3tJv45qUuqSvNKb3vJcz11Itau7bRbhbWys7aS4aEtCixKCrl1hDOygeXE
FkIPQvkxock06WGpyXO0oxT3stuV7ef6PUKuOxF3B1aknJbOpN3fMn72u17PXql1O5t4I7WN
YYVWOONQqoihUUAYAVRwoHYDgVzpKKtFWS2S0t6CnOVSTqVZOU5NuUpNuUm9227tt9W2VrG7
N2ZuAFimaJSO4VVyT77iw49K1lHk5fON/vv+hhGXNfydvy/W4l7pdtqLQvdRiU2somiDZ2rK
FZVfbnazKGYoWB2Mdy4YAiVJxuou11Z+hTina62d16mhUlBQAUAFABQAUAFABQAUAFABQAUA
FABQBn2Gl22meb9ljEZuJXnlOSWklkOWdmYlj/dUZwiBUQKiqopycrXeysvQlRUb2W7u/U0K
koKACgAoAKACgAoAKAMPUP8AQrqG+6I3+jzH0WQgxOfZZfl9hKSeAa3h70ZU+q95fLdfNa/I
wl7soz6fC/ns/v0+ZrzQrOjRSDKOCrD1BGCPyrFPlaa3Rs1dWZ5H9lj067tLN3ezv7abyVuF
Cj7TBLHIkD4YNHKQ3lxyKw8wENtIBBr1+ZzjOaSlCSvy/wAsk05LTVXV2uh51lCUYt8sk7X/
AJk07Ps+ifU6eSfU7LVIjNFHeZtZ1VoGETELLASTHM20HkcLM2ck4GMVypU5U3ytx96Pxara
XVf5G95xmrpS917adV0en4kV3r6Lqdo80F1DtiuQQ0DHk+V0KbwwGDnHTj1pxpP2c1GUXrH7
Xr3sDmueLaktJdPTsP1jxLZyfZgnnErdxHHkTA4Ab1QZPtSp0ZLm2+F/aXl5hOpH3bX+JdH5
i6/rhnsykFrdsWlgwzR+SuftEWPmlK9Tx07/AFopU+WV5SjtLS9/svsOpO8bKMt10t1Xcbrr
aldRQxzmKwiluIgdh82YBGMpYuwWGPaI8k7ZR7iinyRbcbyai99Frptu9/IU+ZpJ2irrzff0
W3mUvDdvb6jqVxd2QL2UBSIXDks11cJuMjb2+Z0hZgu77u8EJwlXVbhCMJ6Td3yrTli9tOjd
vu33JppSm5R+FaX/AJmr3+78zvdQvBYW7zkZKD5VHVnJ2og93cqo9zXDCPPJRWn6Lq/ktTql
Lki5dundvZfNjNLszY2yQscuAWkPrI5LyH6F2bHtinOXNJyW3TyS0X4ChHkio9evq9X+JoVm
aBQBw+q61qF3qn9haL5EUsMC3F3dXCPKkKyMywxpCkkRklkKO3zSoiIuTuLAV0RhGMfaVL2b
sktL23d9bJem5hKUnL2cLKyu29bX2001fqWF1m58O2zP4jlgdjKIrdrOKffc7lBVFtczy+eS
HykTSLtG/KgMFXKpu1FPa75mrL56K3rYfM4L941vpZPX5au/oKfHWjR2hv5Z2hiSdLaRZYZk
lincgLFLC0YliY5By6Ku0hs7eaPZTvypa2urNWaXVO9mHtYW5m7K9tmmn2a3RRb4laIiyFnu
Fe3yZoTZ3YnhQKH86aDyfNig2EN5zqIyDw2ciq9hPTRa7PmjZvsnezfkT7aGu+m65XdebVr2
8zQ1DxvpOmyRwvLJNNcW63UMdvBPcPJAxwJUEMb5XueeF+Y4BBMRpTldpWSdm20rPtqynUjG
yvq1dJJvTvoQ2Pj/AETUpoIbWdpBeELBMIZxbySFC/ki4MYhE+0EmEuJFIKMokG2m6M4ptrb
dXV0u9r3t5iVWDaSe+zs7el9r+W5pN4p0xLGTVTNizt5Hhkk8uX5ZI5vs7rs2bziX5MqpU/e
BK/NU+zlzKFveaulp2v+RfPHlc76LTr0dvzM7U/HmkaTPPazSTPNY7TcrDa3M3kK8ayiSVoo
mVY/LZWMmdo5XO5WAqNGckpJKz2u0r62srvcl1YxbTvdb2Tdr662RaHiO3F88ZubcWsenx3x
+WQMsbySj7Q05P2cwFE+VR+8UqzsdjLS5HyrR35nHpuraW3v+A+dXtdW5eb5a632sVLXx5pV
2jyIblUjhNwrPZXiCWEMieZBugBnG6RABFuY7gQuOabozVlpvb4o6PXR66bdRKrF7X2v8Mld
eWmvyK9x4/sFsr24gE63Gn25uGtri1uYJtpDCJvKkiWRoncbTIisqDJcqATTVGV4p2tJ2umm
vPVO1/Il1Y2k1e6V7NNPy0tsRaP42i1saa0LrC1+WWWKa2u0d5FtDcMls7pGm1CNxlbfFJGp
WNvMIpypOHPf7OzTjp71tV+m/cI1FLltpfo010vpt9+xpQeONJuLpbOOV8ySmCOYwTC1lnUk
GGK6MYt5JMgqFWQ7mBVctxUOlNLmtsr2urpd3G90vkUqkW+VPrZOzs32T2K0vxD0SGR4jNIR
BcNazyrbXJggnWTyik8/leVFmT5VZ3CtwwOwhjSoztey1V0rq7Vr6K92L2sFpfZ2ejsntq7W
WojePbJL02fkXphSbyHvVt2Nkku7YUabORiUiIts2ByMts+cNUZOKleKbV1G/vNb3S9NTleL
hGo6bjUspcrnyP2altZy6Wem1r+Wp3Fcx6IdKACgAoAKADpQAUAV7m2ju4nglG6ORSrD2Iwf
x9D2pxbg1KOjTuiWlJOL2ZlaTdujNp12c3MAyGP/AC3hzhZh6n+GUfwyezLnepFfxYfC+n8s
usf1Xl6MyhJr93P4l/5Muj/z8xde0OHXbZreT5HKkJJjJUn24yMgEjIPAIIYAhUqjpSUlt1X
9f13KqQVRcr+T7Hnt/ez6BNaSXczW0sTmJvtAaW0dZlCM8Vx8siqHEbmOaTKLnC4XnvjFVVN
QV01f3dJprWzjttdXS1+Zxyk6bi5OzTtrrHXs9100b0Ohu7y/wDttjcGGGZd00YaCcFWLwlg
P3ioB/q+OTngZrnjGHJON2tn70ez8m+5s3Lmi7J7rR915+hNrF/evLZx/Y3U/agwHnQ87I5G
I4Y9uefT1pU4xSm+dfD2fVoc5SvFcv2u67MzPE2qXSm2t7v7JYI84lLSzGQqkAMhYoBGpG4K
oAkyWIArSjCPvShzSajayVtZab6/kRUk/dUuWOt9XfRa7afmRW+nT+KLtbiZpZrKFf3csyCK
N5GJy9va7QflT5Uln38sWXdgU3JUIuMUlN7pO7S7Slfvuo28xKLqu7u4rZvTXyj+rPSLa2jt
I1hhUJGgwqjoB/iepPUkknmvObcnd7nakoqy2RhQv/bd0Jl5s7Nj5Z7TTjKlx6xw8qp6NIWI
zsBrpa9jHl+3Jar+WPb1lu/L1Zzr95K6+CL085d/Rfn6HSVynSFABQB5vf8A2nwxr02ri3nu
7DU7aCGY2sbTzQT2rTGNmhQGRoZI5mXdGrlXX5lAYGupWqU1TulKLbV3ZNO19drprqczvTm5
2bjJJO2rTV+nbUo6rfXOo3en6/HY3otdLuLhZIngIuXjuLYxi5itcmYiJyEKFBOVaQrHgENc
YqKlS5o3klZ30Vneze2vrYmTbcaijK0W9La6rdLfT7zAvdLvtYvpdZhtbiKC61fQjHHLE0cx
isZT591JCRviT95tHmBX8uIMwUbRWilGEVTbV1Cps9LyWiT6/LuZuLk3NJpOdPS1naL1dun/
AADrDpt1/auvzeU/l3VhZRwNtOJXSK9Dqh/iZS6AgdCw9aw5koUlfaUr+V3E2s+ao7aOMbee
kjN8G6ReWV/pslxDJEkPhm0tpGZSAk6SRloWJ6SKASV6jFXVknGaTWtWTXo76kU4uLjdWtTS
9H2MzT9Ev4tA0K2aCVZrXV4ppkKHdHGLi5Yu46qoVlJJ4ww9atyj7So01ZwaXm7IlRahTVnd
TTa8rsydQhv4NB1Dw4thfS3j388qtHAxt2hl1AXKSrOcRuDG2DGhaYMDujADMLjyupGrzRUe
VK19bqNrW3X5eZDTUJUuWV+ZvbSzle9/6Z3dvpt0l54kcxOFvPI+znacS7dNiiPln+LEgKHG
fmBHWuZyVqSvte/l77f5HQotOrpva3n7qR5/J4R1S/sfskcDpK3hTS7UCQFFNzBNJJJasxwF
cqAjqxGA43cE11KpGMua+ntpv5NWT/rsc/s5NcqX/LqC+abuv67nba14o1DU9Mlj0az1K0u0
SJ5Ge0KPHH50Szx23nDy57kQtK0XlCRDsO1t5jVueFOMZL2kota297fR2btsr2vf/M2lOUot
QjJPTpa2qva+7te1v8jmbLQ7i91C/ks4tUeG50Ke2jm1MzBpLh5ThFWchoVwR8hjiB+ZwpB3
tq5KMYpuF1UTtC2it5b/AImSi3KTSlZwavK+9/Pb8P1NHTornVT4dCW15bf2aJoLlpreWEwv
/ZUkO75wu5PNYIsikoz8KxqXaHtdYvms1Zp399P8uhavL2dk1y3Tumre41+ZnwWd7PoNl4PF
lcw31rNZpLOYWW1jS0uY5nuo7rAifzUjJRI2MxaTayghqtuKqSr8ycWpWV/efMrWa30v6aEp
PkjR5WmmtbaKzve+2v36lu/0S/fwrr1mkEpuLq/1OSGIId8qS3ZeNkXqyuvzKR1HIqVKKq0p
XVlGF32tHUbi/Z1IpO7lOy73ZR1OwuLbVLg6Taazp2oyzMytaskmlXD7maO4uWkwmHVsyx4A
j5UAvndpBpwiqkqcoJbS0nHvGNu3R9fQ8mrGUa03QhXhUcm1KLvRm7tqdS7tqn70dltq7t+9
jpz1ryz6QKACgAoAKACgAoAKAM7UNOS/VTuMU0R3RTJjfG3TIzwVYcOjZV14I6EaQm6d+sXu
ns1+nk90ZygpeTWzW6f9brqUrbVmgcWupKIJydqOP9TN6eWx+65/55OdwP3d45rSVO656Wse
q+1H1XbzWnoQp8r5Kmj6P7MvR9/J6+pR17XYLVJ7OSPfN5aiGKRAUuXlyqrGDkPtbAlGMqpy
eOaulScnGado3fM07OKWt3202JqVFG8GtbaJ/av27+Zz2paBpNolsZV8tmLO8ls5jRDBE8sk
iqNwCjaV2IBncFreFSpJyttslJXb5mkl0+9mMoQio3++LtaybbIzowuNk8sOoBFSSSIm4Tk+
WSBKoJKF1+VeDhjhuafPy3ipU73Sfuvv072Dlvq4ztZtart17XMvTLSO5dZ9MgtZbiWAusw3
ztAyjzY1kllURfvW/dMsaq6Ft4ztzW03yrlqykoqVraR5r6NpJ30Wqvo9jKKvrTUbtb6u3VX
b01209TvrLxTb3qJLGrrDs3zSuPLjgOOY3Z9u6QN8hVN2DnJFefKhKDcXa97RS1cvNJdLa6n
ZGrGSv0tq3ol5O/X0HM02vfIge3sP4nOUluB/dQcNFER95ziRwcIFB3U/doauzqdFuo+vRvy
2XXsLWrorxh32cvTsvPd9O50MUSQIscahEQBVVRgADgAAcAAVzNtu73OhJJWWiRJSGFABQAU
AFABQAUAFABQAUAFABQAUAFABQAUAFABQAUAFABQAUAFABQAUAFABQBDPbxXKGKZFkjbgq4D
KR7g8U03F3i7NdVoJpSVmrrszCbRrizwdOuCir0huAZoh7IxImjHsHZR0CgV0e0jL+LG/wDe
j7r+f2X9y9TD2bj/AA5WXaXvL5dV9/yMWLRJYHcS2MciukqYiun8tVm5lEcUoAiMh+9sxjtj
Jzu6iaXLUas09YK/u7Xa3t5mKg1e8E9GtJOyvvZPa5NbWWoQvGZFupkt/wDVxvcW6rwpUeYY
1V5doPG7jPLBmwalyg00nFN7tRlf5Xdl8vvKSmrXUmlsnKK++2/9XLNhaanbQJaWyQWcMQCK
ZHa4kCj2URITjplqmUqTbnJyk3rolFfq/wABxVRJQioxS0V25P8ARfiaUGhxh1mvHe8mQ5Vp
cbEPrHCoEaH/AGtpk9XNZuq7ctNKEey3frLd+m3kaKmlrNuTXfZei2X5+ZuVzm4UAFABQAUA
FABQAUAFABQAUAFABQAUAFABQAUAFABQAUAFABQAUAFABQAUAFAH/9k=

--=_reb-r518C6130-t4DD28338--

